library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

package the_snake_game_package is

-- VGA 640-by-480 sync parameters
   	constant HORIZONTAL_DISPLAY: integer:=640; --horizontal display area
   	constant HORIZONTAL_FRONT_PORCH: integer:=16 ; --h. front porch
   	constant HORIZONTAL_BACK_PORCH: integer:=48 ; --h. back porch
   	constant HORIZONTAL_RETRACE: integer:=96 ; --h. retrace
   	constant VERTICAL_DISPLAY: integer:=480; --vertical display area
   	constant VERTICAL_FRONT_PORCH: integer:=10;  --v. front porch
	constant VERTICAL_BACK_PORCH: integer:=33;  --v. back porch
	constant VERTICAL_RETRACE: integer:=2;   --v. retrace

-- Snake parameters
	constant BLOCK_SIZE: integer := 16;
	constant LENGTH_MAX: integer := 128;
	constant MAX_X: integer := 640;
	constant MAX_Y: integer := 480;
	constant HEAD_COLOR: std_logic_vector(2 downto 0):="010";
	constant BODY_COLOR: std_logic_vector(2 downto 0):="010";

-- Items parameters
	type color_array is array(1 to 4) of std_logic_vector(2 downto 0);
	type rom_block is array (0 to 15) of std_logic_vector(0 to 15);
	type rom_array is array (1 to 4) of rom_block;
	constant ITEM_COLOR: color_array := ("100", "110", "100", "101");
	
-- Maps parameters
	constant MAX_WALL_BLOCK: integer := 15;
	constant WALL_COLOR: std_logic_vector(2 downto 0):="100";
	constant BORDER_COLOR: std_logic_vector(2 downto 0):="111";

-- ROMS of in-game objects
	constant ITEM_ROM: rom_array :=
		(
		(
		"0000001110000000",
		"0000000110000000",
		"0000000010000000",
		"0001110010011100",
		"0011111010111110",
		"0111111111111111",
		"0111111111111111",
		"0111111111111111",
		"0111111111111111",
		"0111111111111111",
		"0111111111111111",
		"0111111111111111",
		"0011111111111110",
		"0001111111111100",
		"0000111111111000",
		"0000000000000000"
		),
		(
		"0000000000111000",
		"0000000001111000",
		"0000000011110000",
		"0000000111100000",
		"0000001111100000",
		"0000011111000000",
		"0000111111000000",
		"0001111110000000",
		"0000111110000000",
		"0000011111000000",
		"0000001111000000",
		"0000000111100000",
		"0000000011100000",
		"0000000001110000",
		"0000000000110000",
		"0000000000010000"
		),
		(
		"0000000000000000",
		"0000000000000000",
		"0000000000111000",
		"0000000000111000",
		"0000000001000000",
		"0000000010000000",
		"0000000100000000",
		"0000011111000000",
		"0000111111100000",
		"0001111111110000",
		"0011111111111000",
		"0011111111111000",
		"0001111111110000",
		"0000111111100000",
		"0000011111000000",
		"0000000000000000"
		),
		(
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0001111101111000",
		"0000111111110000",
		"0000011111100000",
		"0000110000110000",
		"0001100000011000",
		"0011000000001100",
		"1111110000111111",
		"1111110000111111",
		"1111110000111111",
		"1111110000111111",
		"1111110000111111"
		)
	);
	
	constant WALL_ROM: rom_block :=
		(
		"1111111100011111",
		"1111111100000111",
		"1111111100000001",
		"1111111100000000",
		"1111111100000000",
		"1111111100000001",
		"1111111100000111",
		"1111111100011111",
		"1111100011111111",
		"1110000011111111",
		"1000000011111111",
		"0000000011111111",
		"0000000011111111",
		"1000000011111111",
		"1110000011111111",
		"1111100011111111"
		);
	
	constant BORDER_ROM: rom_block :=
		(
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000"
		);

	constant SNAKE_HEAD_ROM: rom_block :=
		(
		"0000000000000000",
		"0000111111110000",
		"0001111111111000",
		"0011111111111100",
		"0110001111000110",
		"0110001111000110",
		"0110001111000110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0011111111111100",
		"0001111111111000",
		"0000111111110000",
		"0000000000000000"
		);

	constant SNAKE_ROM: rom_block :=
		(
		"0000000000000000",
		"0000111111110000",
		"0001111111111000",
		"0011111111111100",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0011111111111100",
		"0111111111111100",
		"0111111111111100",
		"0111111111111100",
		"0011111111111100",
		"0011111111111100",
		"0001111111111000",
		"0000000000000000"
		);

	constant LEVEL_PICKER_ROM: rom_block :=
		(
		"0000000110000000",
		"0000001111000000",
		"0000011111100000",
		"0000111111110000",
		"0001111111111000",
		"0011111111111100",
		"0111111111111110",
		"1111111111111111",
		"1111111111111111",
		"0111111111111110",
		"0011111111111100",
		"0001111111111000",
		"0000111111110000",
		"0000011111100000",
		"0000001111000000",
		"0000000110000000"
		);
		
end package the_snake_game_package;