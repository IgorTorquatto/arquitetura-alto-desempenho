library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

library libs;
	use libs.the_snake_game_package.all;
	
entity stages is
	
	port(
		STAGE_SELECT_FROM_TEXT						: in integer range 1 to 7;
		STAGE_SELECT_FROM_LEVEL						: in integer range 1 to 7;
		STATE										: in std_logic;
		PIXEL_X										: in std_logic_vector (9 downto 0);
    	PIXEL_Y										: in std_logic_vector (9 downto 0);
    	ITEM_X										: in unsigned(9 downto 0);
    	ITEM_Y										: in unsigned(9 downto 0);
    	HEAD_X										: in unsigned(9 downto 0);
    	HEAD_Y										: in unsigned(9 downto 0);
    	ITEM_ON_WALL								: out std_logic;
    	HEAD_ON_WALL								: out std_logic;
    	MAP_ON										: out std_logic;
	 	MAP_RGB										: out std_logic_vector (2 downto 0)
	);
end stages;

architecture arch of stages is
	
	-- Placing items requires 10 bits (to obtain 640 px we need 10 bits)
	type wall_pos is array (0 to MAX_WALL_BLOCK) 	of unsigned(9 downto 0);
	signal wall_x									: wall_pos;
	signal wall_y									: wall_pos;
	signal wall_on_temp_1							: std_logic_vector(0 to MAX_WALL_BLOCK-1);
	signal wall_on_temp_2							: std_logic_vector(0 to MAX_WALL_BLOCK);
	signal wall_on_temp_3							: std_logic_vector(0 to MAX_WALL_BLOCK);
	signal wall_on_temp_4							: std_logic_vector(0 to MAX_WALL_BLOCK-1);
	signal item_on_wall_temp_1						: std_logic_vector(0 to MAX_WALL_BLOCK-1);
	signal item_on_wall_temp_2						: std_logic_vector(0 to MAX_WALL_BLOCK);
	signal head_on_wall_temp_1						: std_logic_vector(0 to MAX_WALL_BLOCK-1);
	signal head_on_wall_temp_2						: std_logic_vector(0 to MAX_WALL_BLOCK);
	signal border_on								: std_logic;
	signal stage_select								: integer range 1 to 7;

	begin
	stage_select <= STAGE_SELECT_FROM_TEXT when STATE='1' else STAGE_SELECT_FROM_LEVEL;
	
	-- show border
	border_on			<= '1' when (0 < unsigned(PIXEL_X) and unsigned(PIXEL_X) < 3)
										or (638 < unsigned(PIXEL_X) and unsigned(PIXEL_X) < 641)
										or (0 < unsigned(PIXEL_Y) and unsigned(PIXEL_Y) < 3)
										or (478 < unsigned(PIXEL_Y) and unsigned(PIXEL_Y) < 481)
										or (79 < unsigned(PIXEL_Y) and unsigned(PIXEL_Y) < 82) 
										else '0';
	-- show map
	MAP_ON 				<= 	wall_on_temp_1(0) or border_on;
	MAP_RGB 			<= 	WALL_COLOR when wall_on_temp_4(0)='1' else
			   				BORDER_COLOR when border_on='1' else
			   				"111";
			   
	a0: for i in 0 to MAX_WALL_BLOCK-2 generate
		wall_on_temp_1(i) <= wall_on_temp_2(i) or wall_on_temp_1(i+1);
	end generate;

	wall_on_temp_1(MAX_WALL_BLOCK-1) <= wall_on_temp_2(MAX_WALL_BLOCK-1) or wall_on_temp_2(MAX_WALL_BLOCK);
	a1: for i in 0 to MAX_WALL_BLOCK generate
		wall_on_temp_2(i) <= '1' when (wall_x(i) <= unsigned(PIXEL_X) 
																	and unsigned(PIXEL_X) < wall_x(i)+ BLOCK_SIZE) 
																	and (wall_y(i) <= unsigned(PIXEL_Y) 
																	and unsigned(PIXEL_Y) < wall_y(i)+ BLOCK_SIZE) 
																	else '0';
	end generate;
	
	a3: for i in 0 to MAX_WALL_BLOCK generate
		wall_on_temp_3(i) <= WALL_ROM(to_integer(unsigned(PIXEL_Y(3 downto 0)) - wall_y(i)(3 downto 0)))(to_integer(unsigned(PIXEL_X(3 downto 0)) - wall_x(i)(3 downto 0)));
	end generate;
	
	a4: for i in 0 to MAX_WALL_BLOCK-2 generate
		wall_on_temp_4(i) <= wall_on_temp_3(i) or wall_on_temp_4(i+1);
	end generate;

	wall_on_temp_4(MAX_WALL_BLOCK-1) <= wall_on_temp_3(MAX_WALL_BLOCK-1) or wall_on_temp_3(MAX_WALL_BLOCK);
	
	-- item on wall check
	ITEM_ON_WALL <= item_on_wall_temp_1(0);
	
	b0: for i in 0 to MAX_WALL_BLOCK-2 generate
		item_on_wall_temp_1(i) <= item_on_wall_temp_2(i) or item_on_wall_temp_1(i+1);
	end generate;
	
	item_on_wall_temp_1(MAX_WALL_BLOCK-1) <= item_on_wall_temp_2(MAX_WALL_BLOCK-1) or item_on_wall_temp_2(MAX_WALL_BLOCK);
	b1: for i in 0 to MAX_WALL_BLOCK generate
		item_on_wall_temp_2(i) <= '1' when (wall_x(i)=ITEM_X) and (wall_y(i)=ITEM_Y) else '0';
	end generate;
	
	-- head on wall check
	HEAD_ON_WALL <= head_on_wall_temp_1(0);
	c0: for i in 0 to MAX_WALL_BLOCK-2 generate
		head_on_wall_temp_1(i) <= head_on_wall_temp_2(i) or head_on_wall_temp_1(i+1);
	end generate;
	
	head_on_wall_temp_1(MAX_WALL_BLOCK-1) <= head_on_wall_temp_2(MAX_WALL_BLOCK-1) or head_on_wall_temp_2(MAX_WALL_BLOCK);
	
	c1: for i in 0 to MAX_WALL_BLOCK generate
		head_on_wall_temp_2(i) <= '1' when (wall_x(i)=HEAD_X) and (wall_y(i)=HEAD_Y) else '0';
	end generate;

------------------------------------------------------------------------------------------------------------------------------
-- LEVEL SET 3
	-- Wall Placement on Stage, specify stage as well.
	wall_x(0) <= to_unsigned(272,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
				 
	wall_y(0) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(1) <= to_unsigned(368,10) when stage_select=1 else
				 to_unsigned(1000,10) when stage_select=2 else
				 to_unsigned(0,10);	 
		
	wall_y(1) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(2) <= to_unsigned(416,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
				 
	wall_y(2) <= to_unsigned(192,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(3) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(3) <= to_unsigned(192,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(4) <= to_unsigned(320,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);	 
	
	wall_y(4) <= to_unsigned(192,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(5) <= to_unsigned(272,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);	 
	
	wall_y(5) <= to_unsigned(288,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(6) <= to_unsigned(240,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
				 
	wall_y(6) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(7) <= to_unsigned(240,10) when stage_select=1 else
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(7) <= to_unsigned(256,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(8) <= to_unsigned(240,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(8) <= to_unsigned(288,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(9) <= to_unsigned(320,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(9) <= to_unsigned(320,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(10) <= to_unsigned(400,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(10) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(11) <= to_unsigned(400,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
		
	wall_y(11) <= to_unsigned(288,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------			 
	wall_x(12) <= to_unsigned(416,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else  
				 to_unsigned(0,10);
	
	wall_y(12) <= to_unsigned(320,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------		 
	wall_x(13) <= to_unsigned(400,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
		
	wall_y(13) <= to_unsigned(256,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(14) <= to_unsigned(368,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	
	wall_y(14) <= to_unsigned(288,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
	----------------------------------------------------
	wall_x(15) <= to_unsigned(224,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);
				 
	wall_y(15) <= to_unsigned(320,10) when stage_select=1 else 
				 to_unsigned(1000,10) when stage_select=2 else 
				 to_unsigned(0,10);

end;
